
module niosLab2 (
	buts_export,
	clk_clk,
	leds_name,
	reset_reset_n);	

	input	[3:0]	buts_export;
	input		clk_clk;
	output	[3:0]	leds_name;
	input		reset_reset_n;
endmodule
